hany@hany-Inspiron-3542.5309:1498537505